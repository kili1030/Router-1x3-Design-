package router_pkg;

  import uvm_pkg::*;

	
`include "uvm_macros.svh"
`include "src_agent_config.sv"
`include "dst_agent_config.sv"
`include "env_config.sv"



`include "src_xtn.sv"



`include "src_driver.sv"
`include "src_monitor.sv"
`include "src_sequencer.sv"
`include "src_agent.sv"	
`include "src_agent_top.sv"
`include "src_seqs.sv"

`include "dst_xtn.sv"

`include "dst_driver.sv"	
`include "dst_monitor.sv"	
`include "dst_sequencer.sv"
`include "dst_seqs.sv"	
`include "dst_agent.sv"	
`include "dst_agent_top.sv"

`include "virtual_sequencer.sv"
`include "virtual_seqs.sv"
`include "router_score.sv"	
	

`include "router_env.sv"
`include "router_base_test.sv"			
	

endpackage
